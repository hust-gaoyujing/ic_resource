library verilog;
use verilog.vl_types.all;
entity txblock_tb is
end txblock_tb;
