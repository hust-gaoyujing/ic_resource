library verilog;
use verilog.vl_types.all;
entity rxblock_tb is
end rxblock_tb;
