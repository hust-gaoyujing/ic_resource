library verilog;
use verilog.vl_types.all;
entity uart_tb is
end uart_tb;
