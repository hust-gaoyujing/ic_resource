library verilog;
use verilog.vl_types.all;
entity baud_rate_generator_tb is
end baud_rate_generator_tb;
